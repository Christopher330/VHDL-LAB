`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:58:34 07/02/2016 
// Design Name: 
// Module Name:    lab2_fsm1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module lab2_fsm1(
    input read_ins,
    input read_data,
    input write_data,
    input reset,
    input clk,
    output oe,
    output we
    );


endmodule
